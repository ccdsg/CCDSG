module square_LUT(rst_n,
				  clk,
				  work,
				  pixel,
				  pixel_square
					);
					
input        rst_n,clk    ;
input        work         ;
input  [7:0] pixel        ;
output [15:0] pixel_square;

reg    [15:0] pixel_square;

always @(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		pixel_square <= 16'd0;
	end
	else if(work) begin
		case(pixel)
			8'd0  : pixel_square <= 16'd0;
			8'd1  : pixel_square <= 16'd1;
			8'd2  : pixel_square <= 16'd4;
			8'd3  : pixel_square <= 16'd9;
			8'd4  : pixel_square <= 16'd16;
			8'd5  : pixel_square <= 16'd25;
			8'd6  : pixel_square <= 16'd36;
			8'd7  : pixel_square <= 16'd49;
			8'd8  : pixel_square <= 16'd64;
			8'd9  : pixel_square <= 16'd81;
			8'd10 : pixel_square <= 16'd100;
			8'd11 : pixel_square <= 16'd121;
			8'd12 : pixel_square <= 16'd144;
			8'd13 : pixel_square <= 16'd169;
			8'd14 : pixel_square <= 16'd196;
			8'd15 : pixel_square <= 16'd225;
			8'd16 : pixel_square <= 16'd256;
			8'd17 : pixel_square <= 16'd289;
			8'd18 : pixel_square <= 16'd324;
			8'd19 : pixel_square <= 16'd361;
			8'd20 : pixel_square <= 16'd400;
			8'd21 : pixel_square <= 16'd441;
			8'd22 : pixel_square <= 16'd484;
			8'd23 : pixel_square <= 16'd529;
			8'd24 : pixel_square <= 16'd576;
			8'd25 : pixel_square <= 16'd625;
			8'd26 : pixel_square <= 16'd676;
			8'd27 : pixel_square <= 16'd729;
			8'd28 : pixel_square <= 16'd784;
			8'd29 : pixel_square <= 16'd841;
			8'd30 : pixel_square <= 16'd900;
			8'd31 : pixel_square <= 16'd961;
			8'd32 : pixel_square <= 16'd1024 ;
			8'd33 : pixel_square <= 16'd1089 ;
			8'd34 : pixel_square <= 16'd1156 ;
			8'd35 : pixel_square <= 16'd1225 ;
			8'd36 : pixel_square <= 16'd1296 ;
			8'd37 : pixel_square <= 16'd1369 ;
			8'd38 : pixel_square <= 16'd1444 ;
			8'd39 : pixel_square <= 16'd1521 ;
			8'd40 : pixel_square <= 16'd1600 ;
			8'd41 : pixel_square <= 16'd1681 ;
			8'd42 : pixel_square <= 16'd1764 ;
			8'd43 : pixel_square <= 16'd1849 ;
			8'd44 : pixel_square <= 16'd1936 ;
			8'd45 : pixel_square <= 16'd2025 ;
			8'd46 : pixel_square <= 16'd2116 ;
			8'd47 : pixel_square <= 16'd2209 ;
			8'd48 : pixel_square <= 16'd2304 ;
			8'd49 : pixel_square <= 16'd2401 ;
			8'd50 : pixel_square <= 16'd2500 ;
			8'd51 : pixel_square <= 16'd2601 ;
			8'd52 : pixel_square <= 16'd2704 ;
			8'd53 : pixel_square <= 16'd2809 ;
			8'd54 : pixel_square <= 16'd2916 ;
			8'd55 : pixel_square <= 16'd3025 ;
			8'd56 : pixel_square <= 16'd3136 ;
			8'd57 : pixel_square <= 16'd3249 ;
			8'd58 : pixel_square <= 16'd3364 ;
			8'd59 : pixel_square <= 16'd3481 ;
			8'd60 : pixel_square <= 16'd3600 ;
			8'd61 : pixel_square <= 16'd3721 ;
			8'd62 : pixel_square <= 16'd3844 ;
			8'd63 : pixel_square <= 16'd3969 ;
			8'd64 : pixel_square <= 16'd4096 ;
			8'd65 : pixel_square <= 16'd4225 ;
			8'd66 : pixel_square <= 16'd4356 ;
			8'd67 : pixel_square <= 16'd4489 ;
			8'd68 : pixel_square <= 16'd4624 ;
			8'd69 : pixel_square <= 16'd4761 ;
			8'd70 : pixel_square <= 16'd4900 ;
			8'd71 : pixel_square <= 16'd5041 ;
			8'd72 : pixel_square <= 16'd5184 ;
			8'd73 : pixel_square <= 16'd5329 ;
			8'd74 : pixel_square <= 16'd5476 ;
			8'd75 : pixel_square <= 16'd5625 ;
			8'd76 : pixel_square <= 16'd5776 ;
			8'd77 : pixel_square <= 16'd5929 ;
			8'd78 : pixel_square <= 16'd6084 ;
			8'd79 : pixel_square <= 16'd6241 ;
			8'd80 : pixel_square <= 16'd6400 ;
			8'd81 : pixel_square <= 16'd6561 ;
			8'd82 : pixel_square <= 16'd6724 ;
			8'd83 : pixel_square <= 16'd6889 ;
			8'd84 : pixel_square <= 16'd7056 ;
			8'd85 : pixel_square <= 16'd7225 ;
			8'd86 : pixel_square <= 16'd7396 ;
			8'd87 : pixel_square <= 16'd7569 ;
			8'd88 : pixel_square <= 16'd7744 ;
			8'd89 : pixel_square <= 16'd7921 ;
			8'd90 : pixel_square <= 16'd8100 ;
			8'd91 : pixel_square <= 16'd8281 ;
			8'd92 : pixel_square <= 16'd8464 ;
			8'd93 : pixel_square <= 16'd8649 ;
			8'd94 : pixel_square <= 16'd8836 ;
			8'd95 : pixel_square <= 16'd9025 ;
			8'd96 : pixel_square <= 16'd9216 ;
			8'd97 : pixel_square <= 16'd9409 ;
			8'd98 : pixel_square <= 16'd9604 ;
			8'd99 : pixel_square <= 16'd9801 ;
			8'd100: pixel_square <= 16'd10000;
			8'd101: pixel_square <= 16'd10201;
			8'd102: pixel_square <= 16'd10404;
			8'd103: pixel_square <= 16'd10609;
			8'd104: pixel_square <= 16'd10816;
			8'd105: pixel_square <= 16'd11025;
			8'd106: pixel_square <= 16'd11236;
			8'd107: pixel_square <= 16'd11449;
			8'd108: pixel_square <= 16'd11664;
			8'd109: pixel_square <= 16'd11881;
			8'd110: pixel_square <= 16'd12100;
			8'd111: pixel_square <= 16'd12321;
			8'd112: pixel_square <= 16'd12544;
			8'd113: pixel_square <= 16'd12769;
			8'd114: pixel_square <= 16'd12996;
			8'd115: pixel_square <= 16'd13225;
			8'd116: pixel_square <= 16'd13456;
			8'd117: pixel_square <= 16'd13689;
			8'd118: pixel_square <= 16'd13924;
			8'd119: pixel_square <= 16'd14161;
			8'd120: pixel_square <= 16'd14400;
			8'd121: pixel_square <= 16'd14641;
			8'd122: pixel_square <= 16'd14884;
			8'd123: pixel_square <= 16'd15129;
			8'd124: pixel_square <= 16'd15376;
			8'd125: pixel_square <= 16'd15625;
			8'd126: pixel_square <= 16'd15876;
			8'd127: pixel_square <= 16'd16129;
			8'd128: pixel_square <= 16'd16384;
			8'd129: pixel_square <= 16'd16641;
			8'd130: pixel_square <= 16'd16900;
			8'd131: pixel_square <= 16'd17161;
			8'd132: pixel_square <= 16'd17424;
			8'd133: pixel_square <= 16'd17689;
			8'd134: pixel_square <= 16'd17956;
			8'd135: pixel_square <= 16'd18225;
			8'd136: pixel_square <= 16'd18496;
			8'd137: pixel_square <= 16'd18769;
			8'd138: pixel_square <= 16'd19044;
			8'd139: pixel_square <= 16'd19321;
			8'd140: pixel_square <= 16'd19600;
			8'd141: pixel_square <= 16'd19881;
			8'd142: pixel_square <= 16'd20164;
			8'd143: pixel_square <= 16'd20449;
			8'd144: pixel_square <= 16'd20736;
			8'd145: pixel_square <= 16'd21025;
			8'd146: pixel_square <= 16'd21316;
			8'd147: pixel_square <= 16'd21609;
			8'd148: pixel_square <= 16'd21904;
			8'd149: pixel_square <= 16'd22201;
			8'd150: pixel_square <= 16'd22500;
			8'd151: pixel_square <= 16'd22801;
			8'd152: pixel_square <= 16'd23104;
			8'd153: pixel_square <= 16'd23409;
			8'd154: pixel_square <= 16'd23716;
			8'd155: pixel_square <= 16'd24025;
			8'd156: pixel_square <= 16'd24336;
			8'd157: pixel_square <= 16'd24649;
			8'd158: pixel_square <= 16'd24964;
			8'd159: pixel_square <= 16'd25281;
			8'd160: pixel_square <= 16'd25600;
			8'd161: pixel_square <= 16'd25921;
			8'd162: pixel_square <= 16'd26244;
			8'd163: pixel_square <= 16'd26569;
			8'd164: pixel_square <= 16'd26896;
			8'd165: pixel_square <= 16'd27225;
			8'd166: pixel_square <= 16'd27556;
			8'd167: pixel_square <= 16'd27889;
			8'd168: pixel_square <= 16'd28224;
			8'd169: pixel_square <= 16'd28561;
			8'd170: pixel_square <= 16'd28900;
			8'd171: pixel_square <= 16'd29241;
			8'd172: pixel_square <= 16'd29584;
			8'd173: pixel_square <= 16'd29929;
			8'd174: pixel_square <= 16'd30276;
			8'd175: pixel_square <= 16'd30625;
			8'd176: pixel_square <= 16'd30976;
			8'd177: pixel_square <= 16'd31329;
			8'd178: pixel_square <= 16'd31684;
			8'd179: pixel_square <= 16'd32041;
			8'd180: pixel_square <= 16'd32400;
			8'd181: pixel_square <= 16'd32761;
			8'd182: pixel_square <= 16'd33124;
			8'd183: pixel_square <= 16'd33489;
			8'd184: pixel_square <= 16'd33856;
			8'd185: pixel_square <= 16'd34225;
			8'd186: pixel_square <= 16'd34596;
			8'd187: pixel_square <= 16'd34969;
			8'd188: pixel_square <= 16'd35344;
			8'd189: pixel_square <= 16'd35721;
			8'd190: pixel_square <= 16'd36100;
			8'd191: pixel_square <= 16'd36481;
			8'd192: pixel_square <= 16'd36864;
			8'd193: pixel_square <= 16'd37249;
			8'd194: pixel_square <= 16'd37636;
			8'd195: pixel_square <= 16'd38025;
			8'd196: pixel_square <= 16'd38416;
			8'd197: pixel_square <= 16'd38809;
			8'd198: pixel_square <= 16'd39204;
			8'd199: pixel_square <= 16'd39601;
			8'd200: pixel_square <= 16'd40000;
			8'd201: pixel_square <= 16'd40401;
			8'd202: pixel_square <= 16'd40804;
			8'd203: pixel_square <= 16'd41209;
			8'd204: pixel_square <= 16'd41616;
			8'd205: pixel_square <= 16'd42025;
			8'd206: pixel_square <= 16'd42436;
			8'd207: pixel_square <= 16'd42849;
			8'd208: pixel_square <= 16'd43264;
			8'd209: pixel_square <= 16'd43681;
			8'd210: pixel_square <= 16'd44100;
			8'd211: pixel_square <= 16'd44521;
			8'd212: pixel_square <= 16'd44944;
			8'd213: pixel_square <= 16'd45369;
			8'd214: pixel_square <= 16'd45796;
			8'd215: pixel_square <= 16'd46225;
			8'd216: pixel_square <= 16'd46656;
			8'd217: pixel_square <= 16'd47089;
			8'd218: pixel_square <= 16'd47524;
			8'd219: pixel_square <= 16'd47961;
			8'd220: pixel_square <= 16'd48400;
			8'd221: pixel_square <= 16'd48841;
			8'd222: pixel_square <= 16'd49284;
			8'd223: pixel_square <= 16'd49729;
			8'd224: pixel_square <= 16'd50176;
			8'd225: pixel_square <= 16'd50625;
			8'd226: pixel_square <= 16'd51076;
			8'd227: pixel_square <= 16'd51529;
			8'd228: pixel_square <= 16'd51984;
			8'd229: pixel_square <= 16'd52441;
			8'd230: pixel_square <= 16'd52900;
			8'd231: pixel_square <= 16'd53361;
			8'd232: pixel_square <= 16'd53824;
			8'd233: pixel_square <= 16'd54289;
			8'd234: pixel_square <= 16'd54756;
			8'd235: pixel_square <= 16'd55225;
			8'd236: pixel_square <= 16'd55696;
			8'd237: pixel_square <= 16'd56169;
			8'd238: pixel_square <= 16'd56644;
			8'd239: pixel_square <= 16'd57121;
			8'd240: pixel_square <= 16'd57600;
			8'd241: pixel_square <= 16'd58081;
			8'd242: pixel_square <= 16'd58564;
			8'd243: pixel_square <= 16'd59049;
			8'd244: pixel_square <= 16'd59536;
			8'd245: pixel_square <= 16'd60025;
			8'd246: pixel_square <= 16'd60516;
			8'd247: pixel_square <= 16'd61009;
			8'd248: pixel_square <= 16'd61504;
			8'd249: pixel_square <= 16'd62001;
			8'd250: pixel_square <= 16'd62500;
			8'd251: pixel_square <= 16'd63001;
			8'd252: pixel_square <= 16'd63504;
			8'd253: pixel_square <= 16'd64009;
			8'd254: pixel_square <= 16'd64516;
			8'd255: pixel_square <= 16'd65025;
			default:pixel_square <= 16'd0;
		endcase
	end
	else 
		pixel_square <= 0;
end

endmodule